LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE work.parameters.ALL;

ENTITY testset_demo IS
  PORT (p_pid_out       : OUT REAL RANGE -1.0 TO 1.0;
        t_pid_out       : OUT REAL RANGE -1.0 TO 1.0;
        p_enable    : OUT std_logic;
        t_enable    : OUT std_logic;
        rst       : OUT std_logic;
        clk       : OUT std_logic);
END testset_demo;

ARCHITECTURE set1 OF testset_demo IS
   CONSTANT period_clk : time := 20 ns;
BEGIN
  
  rst <= '1', '0' after 50 ns;
  
  --p_pid_out <= 0.2, -0.6 after 200 ms, 1.0 after 400 ms;
  --t_pid_out <= -0.1, 0.8 after 150 ms, -0.3 after 300 ms;

  p_enable <= '1';
  t_enable <= '1';

  clock_process : PROCESS
   BEGIN
      clk <= '0';
      WAIT FOR period_clk /2;
      clk <= '1';
      WAIT FOR period_clk /2;
   END PROCESS;
   
   t_pid_out <= 0.0,
-0.17	after	30.0	ms,
-0.07	after	40.0	ms,
-0.05	after	50.0	ms,
0.06	after	60.0	ms,
0.00	after	70.0	ms,
0.11	after	80.0	ms,
0.05	after	90.0	ms,
0.06	after	100.0	ms,
0.08	after	110.0	ms,
0.10	after	120.0	ms,
0.02	after	130.0	ms,
0.02	after	140.0	ms,
0.02	after	150.0	ms,
0.02	after	160.0	ms,
0.02	after	170.0	ms,
-0.08	after	180.0	ms,
0.00	after	190.0	ms,
0.00	after	200.0	ms,
0.48	after	210.0	ms,
0.08	after	220.0	ms,
-0.11	after	230.0	ms,
-0.14	after	240.0	ms,
-0.18	after	250.0	ms,
-0.11	after	260.0	ms,
-0.13	after	270.0	ms,
-0.05	after	280.0	ms,
-0.05	after	290.0	ms,
0.05	after	300.0	ms,
0.06	after	310.0	ms,
-0.02	after	320.0	ms,
0.08	after	330.0	ms,
0.00	after	340.0	ms,
0.00	after	350.0	ms,
0.00	after	360.0	ms,
0.09	after	370.0	ms,
0.49	after	380.0	ms,
0.10	after	390.0	ms,
-0.19	after	400.0	ms,
-0.14	after	410.0	ms,
-0.18	after	420.0	ms,
-0.11	after	430.0	ms,
-0.13	after	440.0	ms,
0.43	after	450.0	ms,
0.03	after	460.0	ms,
-0.06	after	470.0	ms,
-0.08	after	480.0	ms,
-0.10	after	490.0	ms,
-0.11	after	500.0	ms,
-0.13	after	510.0	ms,
-0.05	after	520.0	ms,
0.05	after	530.0	ms,
0.54	after	540.0	ms,
0.07	after	550.0	ms,
-0.13	after	560.0	ms,
-0.06	after	570.0	ms,
-0.18	after	580.0	ms,
-0.11	after	590.0	ms,
-0.03	after	600.0	ms,
-0.03	after	610.0	ms,
-0.03	after	620.0	ms,
0.45	after	630.0	ms,
0.05	after	640.0	ms,
-0.05	after	650.0	ms,
-0.06	after	660.0	ms,
-0.18	after	670.0	ms,
-0.11	after	680.0	ms,
-0.03	after	690.0	ms,
-0.03	after	700.0	ms,
-0.03	after	710.0	ms,
-0.03	after	720.0	ms,
0.06	after	730.0	ms,
0.46	after	740.0	ms,
0.07	after	750.0	ms,
-0.03	after	760.0	ms,
-0.14	after	770.0	ms,
-0.08	after	780.0	ms,
-0.10	after	790.0	ms,
-0.11	after	800.0	ms,
-0.13	after	810.0	ms,
-0.05	after	820.0	ms,
0.52	after	830.0	ms,
0.15	after	840.0	ms,
-0.03	after	850.0	ms,
-0.14	after	860.0	ms,
-0.18	after	870.0	ms,
-0.11	after	880.0	ms,
-0.13	after	890.0	ms,
-0.05	after	900.0	ms,
0.05	after	910.0	ms,
-0.03	after	920.0	ms,
0.06	after	930.0	ms,
0.08	after	940.0	ms,
0.48	after	950.0	ms,
0.08	after	960.0	ms,
-0.11	after	970.0	ms,
-0.14	after	980.0	ms,
-0.18	after	990.0	ms,
-0.11	after	1000.0	ms,
-0.03	after	1010.0	ms,
-0.03	after	1020.0	ms,
-0.03	after	1030.0	ms,
-0.03	after	1040.0	ms,
0.06	after	1050.0	ms,
-0.02	after	1060.0	ms,
-0.02	after	1070.0	ms,
0.08	after	1080.0	ms,
0.00	after	1090.0	ms,
0.00	after	1100.0	ms,
0.00	after	1110.0	ms,
0.00	after	1120.0	ms,
0.57	after	1130.0	ms,
0.10	after	1140.0	ms,
-0.10	after	1150.0	ms,
-0.22	after	1160.0	ms,
-0.18	after	1170.0	ms,
-0.11	after	1180.0	ms,
-0.13	after	1190.0	ms,
-0.05	after	1200.0	ms,
-0.05	after	1210.0	ms,
0.05	after	1220.0	ms,
0.06	after	1230.0	ms,
-0.02	after	1240.0	ms,
-0.02	after	1250.0	ms,
0.08	after	1260.0	ms,
0.00	after	1270.0	ms,
0.00	after	1280.0	ms,
0.09	after	1290.0	ms,
0.02	after	1300.0	ms,
0.02	after	1310.0	ms,
-0.08	after	1320.0	ms,
0.00	after	1330.0	ms,
0.00	after	1340.0	ms,
0.00	after	1350.0	ms,
0.00	after	1360.0	ms;
   
   p_pid_out <= 0.0,
0.99	after	30	ms,
0.99	after	40	ms,
0.99	after	50	ms,
0.99	after	60	ms,
0.99	after	70	ms,
0.92	after	80	ms,
0.82	after	90	ms,
0.84	after	100	ms,
0.74	after	110	ms,
0.59	after	120	ms,
0.56	after	130	ms,
0.52	after	140	ms,
0.47	after	150	ms,
0.34	after	160	ms,
0.32	after	170	ms,
0.29	after	180	ms,
0.24	after	190	ms,
0.19	after	200	ms,
0.14	after	210	ms,
0.09	after	220	ms,
0.12	after	230	ms,
0.04	after	240	ms,
0.06	after	250	ms,
0.05	after	260	ms,
-0.05	after	270	ms,
-0.04	after	280	ms,
-0.05	after	290	ms,
-0.07	after	300	ms,
-0.09	after	310	ms,
-0.03	after	320	ms,
-0.09	after	330	ms,
-0.04	after	340	ms,
-0.11	after	350	ms,
-0.07	after	360	ms,
-0.13	after	370	ms,
-0.09	after	380	ms,
-0.07	after	390	ms,
-0.07	after	400	ms,
-0.06	after	410	ms,
-0.06	after	420	ms,
-0.06	after	430	ms,
-0.06	after	440	ms,
-0.06	after	450	ms,
-0.06	after	460	ms,
-0.06	after	470	ms,
-0.06	after	480	ms,
-0.06	after	490	ms,
-0.06	after	500	ms,
-0.06	after	510	ms,
-0.06	after	520	ms,
-0.06	after	530	ms,
-0.06	after	540	ms,
-0.48	after	550	ms,
-0.24	after	560	ms,
-0.2	after	570	ms,
-0.18	after	580	ms,
-0.51	after	590	ms,
-0.8	after	600	ms,
-0.5	after	610	ms,
-0.35	after	620	ms,
-0.69	after	630	ms,
-0.48	after	640	ms,
-0.79	after	650	ms,
-0.57	after	660	ms,
-0.45	after	670	ms,
-0.72	after	680	ms,
-0.55	after	690	ms,
-0.8	after	700	ms,
-0.53	after	710	ms,
-0.89	after	720	ms,
-0.6	after	730	ms,
-0.86	after	740	ms,
-0.61	after	750	ms,
-0.46	after	760	ms,
-0.7	after	770	ms,
-0.5	after	780	ms,
-0.81	after	790	ms,
-0.57	after	800	ms,
-0.43	after	810	ms,
-0.68	after	820	ms,
-0.48	after	830	ms,
-0.36	after	840	ms,
-0.62	after	850	ms,
-0.43	after	860	ms,
-0.73	after	870	ms,
-0.49	after	880	ms,
-0.78	after	890	ms,
-0.11	after	900	ms,
-0.46	after	910	ms,
-0.31	after	920	ms,
-0.64	after	930	ms,
-0.41	after	940	ms,
-0.7	after	950	ms,
-0.45	after	960	ms,
-0.31	after	970	ms,
-0.64	after	980	ms,
-0.41	after	990	ms,
-0.28	after	1000	ms,
-0.19	after	1010	ms,
-0.12	after	1020	ms,
-0.06	after	1030	ms,
-0.01	after	1040	ms,
-0.04	after	1050	ms,
0.05	after	1060	ms,
0.03	after	1070	ms,
0.04	after	1080	ms,
0.05	after	1090	ms,
0.08	after	1100	ms,
0.1	after	1110	ms,
0.13	after	1120	ms,
0.07	after	1130	ms,
0.12	after	1140	ms,
0.08	after	1150	ms,
0.14	after	1160	ms,
0.1	after	1170	ms,
0.09	after	1180	ms,
0.08	after	1190	ms,
0.16	after	1200	ms,
0.12	after	1210	ms,
0.11	after	1220	ms,
0.1	after	1230	ms,
0.1	after	1240	ms,
0.01	after	1250	ms,
0.04	after	1260	ms,
0.06	after	1270	ms,
0.06	after	1280	ms,
0.07	after	1290	ms,
0.07	after	1300	ms,
0.49	after	1310	ms,
-0.09	after	1320	ms,
-0.09	after	1330	ms,
-0.02	after	1340	ms,
0.02	after	1350	ms,
0.03	after	1360	ms,
0.1	after	1370	ms,
0.1	after	1380	ms;

			
END set1;




